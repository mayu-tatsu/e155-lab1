module lab1_mt_testbench();

	logic clk, reset;
	logic [3:0] s;
	logic [2:0] led;
	logic [6:0] seg;
	
endmodule